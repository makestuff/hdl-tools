//
// Copyright (C) 2019 Chris McClelland
//
// Permission is hereby granted, free of charge, to any person obtaining a copy of this software
// and associated documentation files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy, modify, merge, publish,
// distribute, sublicense, and/or sell copies of the Software, and to permit persons to whom the
// Software is furnished to do so, subject to the following conditions:
//
// The above copyright  notice and this permission notice  shall be included in all copies or
// substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR IMPLIED, INCLUDING
// BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM,
// DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.
//
`include "svunit_defines.svh"

`define FATAL_IF(cond, msg) \
  if (cond) begin \
    $display(); \
    $error("\033[31;1mFATAL: %s\033[0m", $sformatf msg); \
    $display(); \
    $stop(1); \
  end

svunit_pkg::svunit_testcase svunit_ut;
localparam string name = NAME;

function void build();
  svunit_ut = new(name);
endfunction

initial begin
  build();
  run();
  $display();
  svunit_ut.report();
  $display();
  if (svunit_ut.get_error_count() > 0) begin
    $error($sformatf("\033[31;1m%0d tests failed\033[0m", svunit_ut.get_error_count()));
    $display();
  end
  $stop();
end
